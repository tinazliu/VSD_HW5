//-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.
//
//
//* File Name : CPU_wrapper.sv
//
//* Purpose :
//
//* Creation Date : 2017-11-05
//
//* Last Modified : Sun 05 Nov 2017 03:45:40 PM CST
//
//* Created By :  Ji-Ying, Li
//
//_._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._
//

`include "AHB_def.svh"

module CPU_wrapper (

);
  
endmodule

