# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : data_array
#       Words            : 64
#       Bits             : 8
#       Byte-Write       : 4
#       Aspect Ratio     : 1
#       Output Loading   : 1.3  (pf)
#       Data Slew        : 2.0  (ns)
#       CK Slew          : 2.0  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2017/10/05 23:56:49
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO data_array
CLASS BLOCK ;
FOREIGN data_array 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 531.960 BY 156.800 ;
SYMMETRY x y r90 ;
#SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 530.840 129.700 531.960 132.940 ;
  LAYER metal3 ;
  RECT 530.840 129.700 531.960 132.940 ;
  LAYER metal2 ;
  RECT 530.840 129.700 531.960 132.940 ;
  LAYER metal1 ;
  RECT 530.840 129.700 531.960 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 121.860 531.960 125.100 ;
  LAYER metal3 ;
  RECT 530.840 121.860 531.960 125.100 ;
  LAYER metal2 ;
  RECT 530.840 121.860 531.960 125.100 ;
  LAYER metal1 ;
  RECT 530.840 121.860 531.960 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 114.020 531.960 117.260 ;
  LAYER metal3 ;
  RECT 530.840 114.020 531.960 117.260 ;
  LAYER metal2 ;
  RECT 530.840 114.020 531.960 117.260 ;
  LAYER metal1 ;
  RECT 530.840 114.020 531.960 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 106.180 531.960 109.420 ;
  LAYER metal3 ;
  RECT 530.840 106.180 531.960 109.420 ;
  LAYER metal2 ;
  RECT 530.840 106.180 531.960 109.420 ;
  LAYER metal1 ;
  RECT 530.840 106.180 531.960 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 98.340 531.960 101.580 ;
  LAYER metal3 ;
  RECT 530.840 98.340 531.960 101.580 ;
  LAYER metal2 ;
  RECT 530.840 98.340 531.960 101.580 ;
  LAYER metal1 ;
  RECT 530.840 98.340 531.960 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 90.500 531.960 93.740 ;
  LAYER metal3 ;
  RECT 530.840 90.500 531.960 93.740 ;
  LAYER metal2 ;
  RECT 530.840 90.500 531.960 93.740 ;
  LAYER metal1 ;
  RECT 530.840 90.500 531.960 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 51.300 531.960 54.540 ;
  LAYER metal3 ;
  RECT 530.840 51.300 531.960 54.540 ;
  LAYER metal2 ;
  RECT 530.840 51.300 531.960 54.540 ;
  LAYER metal1 ;
  RECT 530.840 51.300 531.960 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 43.460 531.960 46.700 ;
  LAYER metal3 ;
  RECT 530.840 43.460 531.960 46.700 ;
  LAYER metal2 ;
  RECT 530.840 43.460 531.960 46.700 ;
  LAYER metal1 ;
  RECT 530.840 43.460 531.960 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 35.620 531.960 38.860 ;
  LAYER metal3 ;
  RECT 530.840 35.620 531.960 38.860 ;
  LAYER metal2 ;
  RECT 530.840 35.620 531.960 38.860 ;
  LAYER metal1 ;
  RECT 530.840 35.620 531.960 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 27.780 531.960 31.020 ;
  LAYER metal3 ;
  RECT 530.840 27.780 531.960 31.020 ;
  LAYER metal2 ;
  RECT 530.840 27.780 531.960 31.020 ;
  LAYER metal1 ;
  RECT 530.840 27.780 531.960 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 19.940 531.960 23.180 ;
  LAYER metal3 ;
  RECT 530.840 19.940 531.960 23.180 ;
  LAYER metal2 ;
  RECT 530.840 19.940 531.960 23.180 ;
  LAYER metal1 ;
  RECT 530.840 19.940 531.960 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 12.100 531.960 15.340 ;
  LAYER metal3 ;
  RECT 530.840 12.100 531.960 15.340 ;
  LAYER metal2 ;
  RECT 530.840 12.100 531.960 15.340 ;
  LAYER metal1 ;
  RECT 530.840 12.100 531.960 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 489.580 155.680 493.120 156.800 ;
  LAYER metal3 ;
  RECT 489.580 155.680 493.120 156.800 ;
  LAYER metal2 ;
  RECT 489.580 155.680 493.120 156.800 ;
  LAYER metal1 ;
  RECT 489.580 155.680 493.120 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 480.900 155.680 484.440 156.800 ;
  LAYER metal3 ;
  RECT 480.900 155.680 484.440 156.800 ;
  LAYER metal2 ;
  RECT 480.900 155.680 484.440 156.800 ;
  LAYER metal1 ;
  RECT 480.900 155.680 484.440 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 472.220 155.680 475.760 156.800 ;
  LAYER metal3 ;
  RECT 472.220 155.680 475.760 156.800 ;
  LAYER metal2 ;
  RECT 472.220 155.680 475.760 156.800 ;
  LAYER metal1 ;
  RECT 472.220 155.680 475.760 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 463.540 155.680 467.080 156.800 ;
  LAYER metal3 ;
  RECT 463.540 155.680 467.080 156.800 ;
  LAYER metal2 ;
  RECT 463.540 155.680 467.080 156.800 ;
  LAYER metal1 ;
  RECT 463.540 155.680 467.080 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 454.860 155.680 458.400 156.800 ;
  LAYER metal3 ;
  RECT 454.860 155.680 458.400 156.800 ;
  LAYER metal2 ;
  RECT 454.860 155.680 458.400 156.800 ;
  LAYER metal1 ;
  RECT 454.860 155.680 458.400 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 446.180 155.680 449.720 156.800 ;
  LAYER metal3 ;
  RECT 446.180 155.680 449.720 156.800 ;
  LAYER metal2 ;
  RECT 446.180 155.680 449.720 156.800 ;
  LAYER metal1 ;
  RECT 446.180 155.680 449.720 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 402.780 155.680 406.320 156.800 ;
  LAYER metal3 ;
  RECT 402.780 155.680 406.320 156.800 ;
  LAYER metal2 ;
  RECT 402.780 155.680 406.320 156.800 ;
  LAYER metal1 ;
  RECT 402.780 155.680 406.320 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 394.100 155.680 397.640 156.800 ;
  LAYER metal3 ;
  RECT 394.100 155.680 397.640 156.800 ;
  LAYER metal2 ;
  RECT 394.100 155.680 397.640 156.800 ;
  LAYER metal1 ;
  RECT 394.100 155.680 397.640 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 385.420 155.680 388.960 156.800 ;
  LAYER metal3 ;
  RECT 385.420 155.680 388.960 156.800 ;
  LAYER metal2 ;
  RECT 385.420 155.680 388.960 156.800 ;
  LAYER metal1 ;
  RECT 385.420 155.680 388.960 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 376.740 155.680 380.280 156.800 ;
  LAYER metal3 ;
  RECT 376.740 155.680 380.280 156.800 ;
  LAYER metal2 ;
  RECT 376.740 155.680 380.280 156.800 ;
  LAYER metal1 ;
  RECT 376.740 155.680 380.280 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 368.060 155.680 371.600 156.800 ;
  LAYER metal3 ;
  RECT 368.060 155.680 371.600 156.800 ;
  LAYER metal2 ;
  RECT 368.060 155.680 371.600 156.800 ;
  LAYER metal1 ;
  RECT 368.060 155.680 371.600 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 359.380 155.680 362.920 156.800 ;
  LAYER metal3 ;
  RECT 359.380 155.680 362.920 156.800 ;
  LAYER metal2 ;
  RECT 359.380 155.680 362.920 156.800 ;
  LAYER metal1 ;
  RECT 359.380 155.680 362.920 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.980 155.680 319.520 156.800 ;
  LAYER metal3 ;
  RECT 315.980 155.680 319.520 156.800 ;
  LAYER metal2 ;
  RECT 315.980 155.680 319.520 156.800 ;
  LAYER metal1 ;
  RECT 315.980 155.680 319.520 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 307.300 155.680 310.840 156.800 ;
  LAYER metal3 ;
  RECT 307.300 155.680 310.840 156.800 ;
  LAYER metal2 ;
  RECT 307.300 155.680 310.840 156.800 ;
  LAYER metal1 ;
  RECT 307.300 155.680 310.840 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 298.620 155.680 302.160 156.800 ;
  LAYER metal3 ;
  RECT 298.620 155.680 302.160 156.800 ;
  LAYER metal2 ;
  RECT 298.620 155.680 302.160 156.800 ;
  LAYER metal1 ;
  RECT 298.620 155.680 302.160 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 289.940 155.680 293.480 156.800 ;
  LAYER metal3 ;
  RECT 289.940 155.680 293.480 156.800 ;
  LAYER metal2 ;
  RECT 289.940 155.680 293.480 156.800 ;
  LAYER metal1 ;
  RECT 289.940 155.680 293.480 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 281.260 155.680 284.800 156.800 ;
  LAYER metal3 ;
  RECT 281.260 155.680 284.800 156.800 ;
  LAYER metal2 ;
  RECT 281.260 155.680 284.800 156.800 ;
  LAYER metal1 ;
  RECT 281.260 155.680 284.800 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 272.580 155.680 276.120 156.800 ;
  LAYER metal3 ;
  RECT 272.580 155.680 276.120 156.800 ;
  LAYER metal2 ;
  RECT 272.580 155.680 276.120 156.800 ;
  LAYER metal1 ;
  RECT 272.580 155.680 276.120 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.180 155.680 232.720 156.800 ;
  LAYER metal3 ;
  RECT 229.180 155.680 232.720 156.800 ;
  LAYER metal2 ;
  RECT 229.180 155.680 232.720 156.800 ;
  LAYER metal1 ;
  RECT 229.180 155.680 232.720 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 220.500 155.680 224.040 156.800 ;
  LAYER metal3 ;
  RECT 220.500 155.680 224.040 156.800 ;
  LAYER metal2 ;
  RECT 220.500 155.680 224.040 156.800 ;
  LAYER metal1 ;
  RECT 220.500 155.680 224.040 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 211.820 155.680 215.360 156.800 ;
  LAYER metal3 ;
  RECT 211.820 155.680 215.360 156.800 ;
  LAYER metal2 ;
  RECT 211.820 155.680 215.360 156.800 ;
  LAYER metal1 ;
  RECT 211.820 155.680 215.360 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 203.140 155.680 206.680 156.800 ;
  LAYER metal3 ;
  RECT 203.140 155.680 206.680 156.800 ;
  LAYER metal2 ;
  RECT 203.140 155.680 206.680 156.800 ;
  LAYER metal1 ;
  RECT 203.140 155.680 206.680 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 194.460 155.680 198.000 156.800 ;
  LAYER metal3 ;
  RECT 194.460 155.680 198.000 156.800 ;
  LAYER metal2 ;
  RECT 194.460 155.680 198.000 156.800 ;
  LAYER metal1 ;
  RECT 194.460 155.680 198.000 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 185.780 155.680 189.320 156.800 ;
  LAYER metal3 ;
  RECT 185.780 155.680 189.320 156.800 ;
  LAYER metal2 ;
  RECT 185.780 155.680 189.320 156.800 ;
  LAYER metal1 ;
  RECT 185.780 155.680 189.320 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 142.380 155.680 145.920 156.800 ;
  LAYER metal3 ;
  RECT 142.380 155.680 145.920 156.800 ;
  LAYER metal2 ;
  RECT 142.380 155.680 145.920 156.800 ;
  LAYER metal1 ;
  RECT 142.380 155.680 145.920 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 133.700 155.680 137.240 156.800 ;
  LAYER metal3 ;
  RECT 133.700 155.680 137.240 156.800 ;
  LAYER metal2 ;
  RECT 133.700 155.680 137.240 156.800 ;
  LAYER metal1 ;
  RECT 133.700 155.680 137.240 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 125.020 155.680 128.560 156.800 ;
  LAYER metal3 ;
  RECT 125.020 155.680 128.560 156.800 ;
  LAYER metal2 ;
  RECT 125.020 155.680 128.560 156.800 ;
  LAYER metal1 ;
  RECT 125.020 155.680 128.560 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 116.340 155.680 119.880 156.800 ;
  LAYER metal3 ;
  RECT 116.340 155.680 119.880 156.800 ;
  LAYER metal2 ;
  RECT 116.340 155.680 119.880 156.800 ;
  LAYER metal1 ;
  RECT 116.340 155.680 119.880 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 107.660 155.680 111.200 156.800 ;
  LAYER metal3 ;
  RECT 107.660 155.680 111.200 156.800 ;
  LAYER metal2 ;
  RECT 107.660 155.680 111.200 156.800 ;
  LAYER metal1 ;
  RECT 107.660 155.680 111.200 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 98.980 155.680 102.520 156.800 ;
  LAYER metal3 ;
  RECT 98.980 155.680 102.520 156.800 ;
  LAYER metal2 ;
  RECT 98.980 155.680 102.520 156.800 ;
  LAYER metal1 ;
  RECT 98.980 155.680 102.520 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 55.580 155.680 59.120 156.800 ;
  LAYER metal3 ;
  RECT 55.580 155.680 59.120 156.800 ;
  LAYER metal2 ;
  RECT 55.580 155.680 59.120 156.800 ;
  LAYER metal1 ;
  RECT 55.580 155.680 59.120 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 46.900 155.680 50.440 156.800 ;
  LAYER metal3 ;
  RECT 46.900 155.680 50.440 156.800 ;
  LAYER metal2 ;
  RECT 46.900 155.680 50.440 156.800 ;
  LAYER metal1 ;
  RECT 46.900 155.680 50.440 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 38.220 155.680 41.760 156.800 ;
  LAYER metal3 ;
  RECT 38.220 155.680 41.760 156.800 ;
  LAYER metal2 ;
  RECT 38.220 155.680 41.760 156.800 ;
  LAYER metal1 ;
  RECT 38.220 155.680 41.760 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 29.540 155.680 33.080 156.800 ;
  LAYER metal3 ;
  RECT 29.540 155.680 33.080 156.800 ;
  LAYER metal2 ;
  RECT 29.540 155.680 33.080 156.800 ;
  LAYER metal1 ;
  RECT 29.540 155.680 33.080 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 20.860 155.680 24.400 156.800 ;
  LAYER metal3 ;
  RECT 20.860 155.680 24.400 156.800 ;
  LAYER metal2 ;
  RECT 20.860 155.680 24.400 156.800 ;
  LAYER metal1 ;
  RECT 20.860 155.680 24.400 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 12.180 155.680 15.720 156.800 ;
  LAYER metal3 ;
  RECT 12.180 155.680 15.720 156.800 ;
  LAYER metal2 ;
  RECT 12.180 155.680 15.720 156.800 ;
  LAYER metal1 ;
  RECT 12.180 155.680 15.720 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 511.900 0.000 515.440 1.120 ;
  LAYER metal3 ;
  RECT 511.900 0.000 515.440 1.120 ;
  LAYER metal2 ;
  RECT 511.900 0.000 515.440 1.120 ;
  LAYER metal1 ;
  RECT 511.900 0.000 515.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 385.420 0.000 388.960 1.120 ;
  LAYER metal3 ;
  RECT 385.420 0.000 388.960 1.120 ;
  LAYER metal2 ;
  RECT 385.420 0.000 388.960 1.120 ;
  LAYER metal1 ;
  RECT 385.420 0.000 388.960 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 369.300 0.000 372.840 1.120 ;
  LAYER metal3 ;
  RECT 369.300 0.000 372.840 1.120 ;
  LAYER metal2 ;
  RECT 369.300 0.000 372.840 1.120 ;
  LAYER metal1 ;
  RECT 369.300 0.000 372.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 342.640 0.000 346.180 1.120 ;
  LAYER metal3 ;
  RECT 342.640 0.000 346.180 1.120 ;
  LAYER metal2 ;
  RECT 342.640 0.000 346.180 1.120 ;
  LAYER metal1 ;
  RECT 342.640 0.000 346.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 320.940 0.000 324.480 1.120 ;
  LAYER metal3 ;
  RECT 320.940 0.000 324.480 1.120 ;
  LAYER metal2 ;
  RECT 320.940 0.000 324.480 1.120 ;
  LAYER metal1 ;
  RECT 320.940 0.000 324.480 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 276.300 0.000 279.840 1.120 ;
  LAYER metal3 ;
  RECT 276.300 0.000 279.840 1.120 ;
  LAYER metal2 ;
  RECT 276.300 0.000 279.840 1.120 ;
  LAYER metal1 ;
  RECT 276.300 0.000 279.840 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 267.620 0.000 271.160 1.120 ;
  LAYER metal3 ;
  RECT 267.620 0.000 271.160 1.120 ;
  LAYER metal2 ;
  RECT 267.620 0.000 271.160 1.120 ;
  LAYER metal1 ;
  RECT 267.620 0.000 271.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 156.640 0.000 160.180 1.120 ;
  LAYER metal3 ;
  RECT 156.640 0.000 160.180 1.120 ;
  LAYER metal2 ;
  RECT 156.640 0.000 160.180 1.120 ;
  LAYER metal1 ;
  RECT 156.640 0.000 160.180 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal3 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal2 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal1 ;
  RECT 139.900 0.000 143.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 530.840 125.780 531.960 129.020 ;
  LAYER metal3 ;
  RECT 530.840 125.780 531.960 129.020 ;
  LAYER metal2 ;
  RECT 530.840 125.780 531.960 129.020 ;
  LAYER metal1 ;
  RECT 530.840 125.780 531.960 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 117.940 531.960 121.180 ;
  LAYER metal3 ;
  RECT 530.840 117.940 531.960 121.180 ;
  LAYER metal2 ;
  RECT 530.840 117.940 531.960 121.180 ;
  LAYER metal1 ;
  RECT 530.840 117.940 531.960 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 110.100 531.960 113.340 ;
  LAYER metal3 ;
  RECT 530.840 110.100 531.960 113.340 ;
  LAYER metal2 ;
  RECT 530.840 110.100 531.960 113.340 ;
  LAYER metal1 ;
  RECT 530.840 110.100 531.960 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 102.260 531.960 105.500 ;
  LAYER metal3 ;
  RECT 530.840 102.260 531.960 105.500 ;
  LAYER metal2 ;
  RECT 530.840 102.260 531.960 105.500 ;
  LAYER metal1 ;
  RECT 530.840 102.260 531.960 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 94.420 531.960 97.660 ;
  LAYER metal3 ;
  RECT 530.840 94.420 531.960 97.660 ;
  LAYER metal2 ;
  RECT 530.840 94.420 531.960 97.660 ;
  LAYER metal1 ;
  RECT 530.840 94.420 531.960 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 86.580 531.960 89.820 ;
  LAYER metal3 ;
  RECT 530.840 86.580 531.960 89.820 ;
  LAYER metal2 ;
  RECT 530.840 86.580 531.960 89.820 ;
  LAYER metal1 ;
  RECT 530.840 86.580 531.960 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 47.380 531.960 50.620 ;
  LAYER metal3 ;
  RECT 530.840 47.380 531.960 50.620 ;
  LAYER metal2 ;
  RECT 530.840 47.380 531.960 50.620 ;
  LAYER metal1 ;
  RECT 530.840 47.380 531.960 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 39.540 531.960 42.780 ;
  LAYER metal3 ;
  RECT 530.840 39.540 531.960 42.780 ;
  LAYER metal2 ;
  RECT 530.840 39.540 531.960 42.780 ;
  LAYER metal1 ;
  RECT 530.840 39.540 531.960 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 31.700 531.960 34.940 ;
  LAYER metal3 ;
  RECT 530.840 31.700 531.960 34.940 ;
  LAYER metal2 ;
  RECT 530.840 31.700 531.960 34.940 ;
  LAYER metal1 ;
  RECT 530.840 31.700 531.960 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 23.860 531.960 27.100 ;
  LAYER metal3 ;
  RECT 530.840 23.860 531.960 27.100 ;
  LAYER metal2 ;
  RECT 530.840 23.860 531.960 27.100 ;
  LAYER metal1 ;
  RECT 530.840 23.860 531.960 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 16.020 531.960 19.260 ;
  LAYER metal3 ;
  RECT 530.840 16.020 531.960 19.260 ;
  LAYER metal2 ;
  RECT 530.840 16.020 531.960 19.260 ;
  LAYER metal1 ;
  RECT 530.840 16.020 531.960 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.840 8.180 531.960 11.420 ;
  LAYER metal3 ;
  RECT 530.840 8.180 531.960 11.420 ;
  LAYER metal2 ;
  RECT 530.840 8.180 531.960 11.420 ;
  LAYER metal1 ;
  RECT 530.840 8.180 531.960 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 485.240 155.680 488.780 156.800 ;
  LAYER metal3 ;
  RECT 485.240 155.680 488.780 156.800 ;
  LAYER metal2 ;
  RECT 485.240 155.680 488.780 156.800 ;
  LAYER metal1 ;
  RECT 485.240 155.680 488.780 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 476.560 155.680 480.100 156.800 ;
  LAYER metal3 ;
  RECT 476.560 155.680 480.100 156.800 ;
  LAYER metal2 ;
  RECT 476.560 155.680 480.100 156.800 ;
  LAYER metal1 ;
  RECT 476.560 155.680 480.100 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 467.880 155.680 471.420 156.800 ;
  LAYER metal3 ;
  RECT 467.880 155.680 471.420 156.800 ;
  LAYER metal2 ;
  RECT 467.880 155.680 471.420 156.800 ;
  LAYER metal1 ;
  RECT 467.880 155.680 471.420 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 459.200 155.680 462.740 156.800 ;
  LAYER metal3 ;
  RECT 459.200 155.680 462.740 156.800 ;
  LAYER metal2 ;
  RECT 459.200 155.680 462.740 156.800 ;
  LAYER metal1 ;
  RECT 459.200 155.680 462.740 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 450.520 155.680 454.060 156.800 ;
  LAYER metal3 ;
  RECT 450.520 155.680 454.060 156.800 ;
  LAYER metal2 ;
  RECT 450.520 155.680 454.060 156.800 ;
  LAYER metal1 ;
  RECT 450.520 155.680 454.060 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 441.840 155.680 445.380 156.800 ;
  LAYER metal3 ;
  RECT 441.840 155.680 445.380 156.800 ;
  LAYER metal2 ;
  RECT 441.840 155.680 445.380 156.800 ;
  LAYER metal1 ;
  RECT 441.840 155.680 445.380 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 398.440 155.680 401.980 156.800 ;
  LAYER metal3 ;
  RECT 398.440 155.680 401.980 156.800 ;
  LAYER metal2 ;
  RECT 398.440 155.680 401.980 156.800 ;
  LAYER metal1 ;
  RECT 398.440 155.680 401.980 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 389.760 155.680 393.300 156.800 ;
  LAYER metal3 ;
  RECT 389.760 155.680 393.300 156.800 ;
  LAYER metal2 ;
  RECT 389.760 155.680 393.300 156.800 ;
  LAYER metal1 ;
  RECT 389.760 155.680 393.300 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 381.080 155.680 384.620 156.800 ;
  LAYER metal3 ;
  RECT 381.080 155.680 384.620 156.800 ;
  LAYER metal2 ;
  RECT 381.080 155.680 384.620 156.800 ;
  LAYER metal1 ;
  RECT 381.080 155.680 384.620 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 372.400 155.680 375.940 156.800 ;
  LAYER metal3 ;
  RECT 372.400 155.680 375.940 156.800 ;
  LAYER metal2 ;
  RECT 372.400 155.680 375.940 156.800 ;
  LAYER metal1 ;
  RECT 372.400 155.680 375.940 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 363.720 155.680 367.260 156.800 ;
  LAYER metal3 ;
  RECT 363.720 155.680 367.260 156.800 ;
  LAYER metal2 ;
  RECT 363.720 155.680 367.260 156.800 ;
  LAYER metal1 ;
  RECT 363.720 155.680 367.260 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 355.040 155.680 358.580 156.800 ;
  LAYER metal3 ;
  RECT 355.040 155.680 358.580 156.800 ;
  LAYER metal2 ;
  RECT 355.040 155.680 358.580 156.800 ;
  LAYER metal1 ;
  RECT 355.040 155.680 358.580 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 311.640 155.680 315.180 156.800 ;
  LAYER metal3 ;
  RECT 311.640 155.680 315.180 156.800 ;
  LAYER metal2 ;
  RECT 311.640 155.680 315.180 156.800 ;
  LAYER metal1 ;
  RECT 311.640 155.680 315.180 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 302.960 155.680 306.500 156.800 ;
  LAYER metal3 ;
  RECT 302.960 155.680 306.500 156.800 ;
  LAYER metal2 ;
  RECT 302.960 155.680 306.500 156.800 ;
  LAYER metal1 ;
  RECT 302.960 155.680 306.500 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 294.280 155.680 297.820 156.800 ;
  LAYER metal3 ;
  RECT 294.280 155.680 297.820 156.800 ;
  LAYER metal2 ;
  RECT 294.280 155.680 297.820 156.800 ;
  LAYER metal1 ;
  RECT 294.280 155.680 297.820 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 285.600 155.680 289.140 156.800 ;
  LAYER metal3 ;
  RECT 285.600 155.680 289.140 156.800 ;
  LAYER metal2 ;
  RECT 285.600 155.680 289.140 156.800 ;
  LAYER metal1 ;
  RECT 285.600 155.680 289.140 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 276.920 155.680 280.460 156.800 ;
  LAYER metal3 ;
  RECT 276.920 155.680 280.460 156.800 ;
  LAYER metal2 ;
  RECT 276.920 155.680 280.460 156.800 ;
  LAYER metal1 ;
  RECT 276.920 155.680 280.460 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 268.240 155.680 271.780 156.800 ;
  LAYER metal3 ;
  RECT 268.240 155.680 271.780 156.800 ;
  LAYER metal2 ;
  RECT 268.240 155.680 271.780 156.800 ;
  LAYER metal1 ;
  RECT 268.240 155.680 271.780 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 224.840 155.680 228.380 156.800 ;
  LAYER metal3 ;
  RECT 224.840 155.680 228.380 156.800 ;
  LAYER metal2 ;
  RECT 224.840 155.680 228.380 156.800 ;
  LAYER metal1 ;
  RECT 224.840 155.680 228.380 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 216.160 155.680 219.700 156.800 ;
  LAYER metal3 ;
  RECT 216.160 155.680 219.700 156.800 ;
  LAYER metal2 ;
  RECT 216.160 155.680 219.700 156.800 ;
  LAYER metal1 ;
  RECT 216.160 155.680 219.700 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 207.480 155.680 211.020 156.800 ;
  LAYER metal3 ;
  RECT 207.480 155.680 211.020 156.800 ;
  LAYER metal2 ;
  RECT 207.480 155.680 211.020 156.800 ;
  LAYER metal1 ;
  RECT 207.480 155.680 211.020 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 198.800 155.680 202.340 156.800 ;
  LAYER metal3 ;
  RECT 198.800 155.680 202.340 156.800 ;
  LAYER metal2 ;
  RECT 198.800 155.680 202.340 156.800 ;
  LAYER metal1 ;
  RECT 198.800 155.680 202.340 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 190.120 155.680 193.660 156.800 ;
  LAYER metal3 ;
  RECT 190.120 155.680 193.660 156.800 ;
  LAYER metal2 ;
  RECT 190.120 155.680 193.660 156.800 ;
  LAYER metal1 ;
  RECT 190.120 155.680 193.660 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 181.440 155.680 184.980 156.800 ;
  LAYER metal3 ;
  RECT 181.440 155.680 184.980 156.800 ;
  LAYER metal2 ;
  RECT 181.440 155.680 184.980 156.800 ;
  LAYER metal1 ;
  RECT 181.440 155.680 184.980 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 138.040 155.680 141.580 156.800 ;
  LAYER metal3 ;
  RECT 138.040 155.680 141.580 156.800 ;
  LAYER metal2 ;
  RECT 138.040 155.680 141.580 156.800 ;
  LAYER metal1 ;
  RECT 138.040 155.680 141.580 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 129.360 155.680 132.900 156.800 ;
  LAYER metal3 ;
  RECT 129.360 155.680 132.900 156.800 ;
  LAYER metal2 ;
  RECT 129.360 155.680 132.900 156.800 ;
  LAYER metal1 ;
  RECT 129.360 155.680 132.900 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 120.680 155.680 124.220 156.800 ;
  LAYER metal3 ;
  RECT 120.680 155.680 124.220 156.800 ;
  LAYER metal2 ;
  RECT 120.680 155.680 124.220 156.800 ;
  LAYER metal1 ;
  RECT 120.680 155.680 124.220 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 112.000 155.680 115.540 156.800 ;
  LAYER metal3 ;
  RECT 112.000 155.680 115.540 156.800 ;
  LAYER metal2 ;
  RECT 112.000 155.680 115.540 156.800 ;
  LAYER metal1 ;
  RECT 112.000 155.680 115.540 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 103.320 155.680 106.860 156.800 ;
  LAYER metal3 ;
  RECT 103.320 155.680 106.860 156.800 ;
  LAYER metal2 ;
  RECT 103.320 155.680 106.860 156.800 ;
  LAYER metal1 ;
  RECT 103.320 155.680 106.860 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 94.640 155.680 98.180 156.800 ;
  LAYER metal3 ;
  RECT 94.640 155.680 98.180 156.800 ;
  LAYER metal2 ;
  RECT 94.640 155.680 98.180 156.800 ;
  LAYER metal1 ;
  RECT 94.640 155.680 98.180 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 51.240 155.680 54.780 156.800 ;
  LAYER metal3 ;
  RECT 51.240 155.680 54.780 156.800 ;
  LAYER metal2 ;
  RECT 51.240 155.680 54.780 156.800 ;
  LAYER metal1 ;
  RECT 51.240 155.680 54.780 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 42.560 155.680 46.100 156.800 ;
  LAYER metal3 ;
  RECT 42.560 155.680 46.100 156.800 ;
  LAYER metal2 ;
  RECT 42.560 155.680 46.100 156.800 ;
  LAYER metal1 ;
  RECT 42.560 155.680 46.100 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 33.880 155.680 37.420 156.800 ;
  LAYER metal3 ;
  RECT 33.880 155.680 37.420 156.800 ;
  LAYER metal2 ;
  RECT 33.880 155.680 37.420 156.800 ;
  LAYER metal1 ;
  RECT 33.880 155.680 37.420 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 25.200 155.680 28.740 156.800 ;
  LAYER metal3 ;
  RECT 25.200 155.680 28.740 156.800 ;
  LAYER metal2 ;
  RECT 25.200 155.680 28.740 156.800 ;
  LAYER metal1 ;
  RECT 25.200 155.680 28.740 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 16.520 155.680 20.060 156.800 ;
  LAYER metal3 ;
  RECT 16.520 155.680 20.060 156.800 ;
  LAYER metal2 ;
  RECT 16.520 155.680 20.060 156.800 ;
  LAYER metal1 ;
  RECT 16.520 155.680 20.060 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 7.840 155.680 11.380 156.800 ;
  LAYER metal3 ;
  RECT 7.840 155.680 11.380 156.800 ;
  LAYER metal2 ;
  RECT 7.840 155.680 11.380 156.800 ;
  LAYER metal1 ;
  RECT 7.840 155.680 11.380 156.800 ;
 END
 PORT
  LAYER metal4 ;
  RECT 520.580 0.000 524.120 1.120 ;
  LAYER metal3 ;
  RECT 520.580 0.000 524.120 1.120 ;
  LAYER metal2 ;
  RECT 520.580 0.000 524.120 1.120 ;
  LAYER metal1 ;
  RECT 520.580 0.000 524.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 498.880 0.000 502.420 1.120 ;
  LAYER metal3 ;
  RECT 498.880 0.000 502.420 1.120 ;
  LAYER metal2 ;
  RECT 498.880 0.000 502.420 1.120 ;
  LAYER metal1 ;
  RECT 498.880 0.000 502.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 377.360 0.000 380.900 1.120 ;
  LAYER metal3 ;
  RECT 377.360 0.000 380.900 1.120 ;
  LAYER metal2 ;
  RECT 377.360 0.000 380.900 1.120 ;
  LAYER metal1 ;
  RECT 377.360 0.000 380.900 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 355.660 0.000 359.200 1.120 ;
  LAYER metal3 ;
  RECT 355.660 0.000 359.200 1.120 ;
  LAYER metal2 ;
  RECT 355.660 0.000 359.200 1.120 ;
  LAYER metal1 ;
  RECT 355.660 0.000 359.200 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 329.000 0.000 332.540 1.120 ;
  LAYER metal3 ;
  RECT 329.000 0.000 332.540 1.120 ;
  LAYER metal2 ;
  RECT 329.000 0.000 332.540 1.120 ;
  LAYER metal1 ;
  RECT 329.000 0.000 332.540 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 312.260 0.000 315.800 1.120 ;
  LAYER metal3 ;
  RECT 312.260 0.000 315.800 1.120 ;
  LAYER metal2 ;
  RECT 312.260 0.000 315.800 1.120 ;
  LAYER metal1 ;
  RECT 312.260 0.000 315.800 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 271.960 0.000 275.500 1.120 ;
  LAYER metal3 ;
  RECT 271.960 0.000 275.500 1.120 ;
  LAYER metal2 ;
  RECT 271.960 0.000 275.500 1.120 ;
  LAYER metal1 ;
  RECT 271.960 0.000 275.500 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 263.280 0.000 266.820 1.120 ;
  LAYER metal3 ;
  RECT 263.280 0.000 266.820 1.120 ;
  LAYER metal2 ;
  RECT 263.280 0.000 266.820 1.120 ;
  LAYER metal1 ;
  RECT 263.280 0.000 266.820 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 148.580 0.000 152.120 1.120 ;
  LAYER metal3 ;
  RECT 148.580 0.000 152.120 1.120 ;
  LAYER metal2 ;
  RECT 148.580 0.000 152.120 1.120 ;
  LAYER metal1 ;
  RECT 148.580 0.000 152.120 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END VCC
PIN DO[31]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 518.380 0.000 519.500 1.120 ;
  LAYER metal3 ;
  RECT 518.380 0.000 519.500 1.120 ;
  LAYER metal2 ;
  RECT 518.380 0.000 519.500 1.120 ;
  LAYER metal1 ;
  RECT 518.380 0.000 519.500 1.120 ;
 END
END DO[31]
PIN DI[31]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER metal3 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER metal2 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER metal1 ;
  RECT 509.700 0.000 510.820 1.120 ;
 END
END DI[31]
PIN DO[30]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 504.740 0.000 505.860 1.120 ;
  LAYER metal3 ;
  RECT 504.740 0.000 505.860 1.120 ;
  LAYER metal2 ;
  RECT 504.740 0.000 505.860 1.120 ;
  LAYER metal1 ;
  RECT 504.740 0.000 505.860 1.120 ;
 END
END DO[30]
PIN DI[30]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER metal3 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER metal2 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER metal1 ;
  RECT 496.680 0.000 497.800 1.120 ;
 END
END DI[30]
PIN DO[29]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER metal3 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER metal2 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER metal1 ;
  RECT 488.000 0.000 489.120 1.120 ;
 END
END DO[29]
PIN DI[29]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 479.940 0.000 481.060 1.120 ;
  LAYER metal3 ;
  RECT 479.940 0.000 481.060 1.120 ;
  LAYER metal2 ;
  RECT 479.940 0.000 481.060 1.120 ;
  LAYER metal1 ;
  RECT 479.940 0.000 481.060 1.120 ;
 END
END DI[29]
PIN DO[28]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 474.980 0.000 476.100 1.120 ;
  LAYER metal3 ;
  RECT 474.980 0.000 476.100 1.120 ;
  LAYER metal2 ;
  RECT 474.980 0.000 476.100 1.120 ;
  LAYER metal1 ;
  RECT 474.980 0.000 476.100 1.120 ;
 END
END DO[28]
PIN DI[28]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 466.300 0.000 467.420 1.120 ;
  LAYER metal3 ;
  RECT 466.300 0.000 467.420 1.120 ;
  LAYER metal2 ;
  RECT 466.300 0.000 467.420 1.120 ;
  LAYER metal1 ;
  RECT 466.300 0.000 467.420 1.120 ;
 END
END DI[28]
PIN DO[27]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 461.960 0.000 463.080 1.120 ;
  LAYER metal3 ;
  RECT 461.960 0.000 463.080 1.120 ;
  LAYER metal2 ;
  RECT 461.960 0.000 463.080 1.120 ;
  LAYER metal1 ;
  RECT 461.960 0.000 463.080 1.120 ;
 END
END DO[27]
PIN DI[27]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 453.280 0.000 454.400 1.120 ;
  LAYER metal3 ;
  RECT 453.280 0.000 454.400 1.120 ;
  LAYER metal2 ;
  RECT 453.280 0.000 454.400 1.120 ;
  LAYER metal1 ;
  RECT 453.280 0.000 454.400 1.120 ;
 END
END DI[27]
PIN DO[26]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 448.320 0.000 449.440 1.120 ;
  LAYER metal3 ;
  RECT 448.320 0.000 449.440 1.120 ;
  LAYER metal2 ;
  RECT 448.320 0.000 449.440 1.120 ;
  LAYER metal1 ;
  RECT 448.320 0.000 449.440 1.120 ;
 END
END DO[26]
PIN DI[26]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 440.260 0.000 441.380 1.120 ;
  LAYER metal3 ;
  RECT 440.260 0.000 441.380 1.120 ;
  LAYER metal2 ;
  RECT 440.260 0.000 441.380 1.120 ;
  LAYER metal1 ;
  RECT 440.260 0.000 441.380 1.120 ;
 END
END DI[26]
PIN DO[25]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 431.580 0.000 432.700 1.120 ;
  LAYER metal3 ;
  RECT 431.580 0.000 432.700 1.120 ;
  LAYER metal2 ;
  RECT 431.580 0.000 432.700 1.120 ;
  LAYER metal1 ;
  RECT 431.580 0.000 432.700 1.120 ;
 END
END DO[25]
PIN DI[25]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 423.520 0.000 424.640 1.120 ;
  LAYER metal3 ;
  RECT 423.520 0.000 424.640 1.120 ;
  LAYER metal2 ;
  RECT 423.520 0.000 424.640 1.120 ;
  LAYER metal1 ;
  RECT 423.520 0.000 424.640 1.120 ;
 END
END DI[25]
PIN DO[24]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 418.560 0.000 419.680 1.120 ;
  LAYER metal3 ;
  RECT 418.560 0.000 419.680 1.120 ;
  LAYER metal2 ;
  RECT 418.560 0.000 419.680 1.120 ;
  LAYER metal1 ;
  RECT 418.560 0.000 419.680 1.120 ;
 END
END DO[24]
PIN WEB[3]
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 414.220 0.000 415.340 1.120 ;
  LAYER metal3 ;
  RECT 414.220 0.000 415.340 1.120 ;
  LAYER metal2 ;
  RECT 414.220 0.000 415.340 1.120 ;
  LAYER metal1 ;
  RECT 414.220 0.000 415.340 1.120 ;
 END
END WEB[3]
PIN DI[24]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 409.880 0.000 411.000 1.120 ;
  LAYER metal3 ;
  RECT 409.880 0.000 411.000 1.120 ;
  LAYER metal2 ;
  RECT 409.880 0.000 411.000 1.120 ;
  LAYER metal1 ;
  RECT 409.880 0.000 411.000 1.120 ;
 END
END DI[24]
PIN DO[23]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 404.920 0.000 406.040 1.120 ;
  LAYER metal3 ;
  RECT 404.920 0.000 406.040 1.120 ;
  LAYER metal2 ;
  RECT 404.920 0.000 406.040 1.120 ;
  LAYER metal1 ;
  RECT 404.920 0.000 406.040 1.120 ;
 END
END DO[23]
PIN DI[23]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 396.860 0.000 397.980 1.120 ;
  LAYER metal3 ;
  RECT 396.860 0.000 397.980 1.120 ;
  LAYER metal2 ;
  RECT 396.860 0.000 397.980 1.120 ;
  LAYER metal1 ;
  RECT 396.860 0.000 397.980 1.120 ;
 END
END DI[23]
PIN DO[22]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 391.900 0.000 393.020 1.120 ;
  LAYER metal3 ;
  RECT 391.900 0.000 393.020 1.120 ;
  LAYER metal2 ;
  RECT 391.900 0.000 393.020 1.120 ;
  LAYER metal1 ;
  RECT 391.900 0.000 393.020 1.120 ;
 END
END DO[22]
PIN DI[22]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 383.220 0.000 384.340 1.120 ;
  LAYER metal3 ;
  RECT 383.220 0.000 384.340 1.120 ;
  LAYER metal2 ;
  RECT 383.220 0.000 384.340 1.120 ;
  LAYER metal1 ;
  RECT 383.220 0.000 384.340 1.120 ;
 END
END DI[22]
PIN DO[21]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 375.160 0.000 376.280 1.120 ;
  LAYER metal3 ;
  RECT 375.160 0.000 376.280 1.120 ;
  LAYER metal2 ;
  RECT 375.160 0.000 376.280 1.120 ;
  LAYER metal1 ;
  RECT 375.160 0.000 376.280 1.120 ;
 END
END DO[21]
PIN DI[21]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 367.100 0.000 368.220 1.120 ;
  LAYER metal3 ;
  RECT 367.100 0.000 368.220 1.120 ;
  LAYER metal2 ;
  RECT 367.100 0.000 368.220 1.120 ;
  LAYER metal1 ;
  RECT 367.100 0.000 368.220 1.120 ;
 END
END DI[21]
PIN DO[20]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal3 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal2 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal1 ;
  RECT 362.140 0.000 363.260 1.120 ;
 END
END DO[20]
PIN DI[20]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 353.460 0.000 354.580 1.120 ;
  LAYER metal3 ;
  RECT 353.460 0.000 354.580 1.120 ;
  LAYER metal2 ;
  RECT 353.460 0.000 354.580 1.120 ;
  LAYER metal1 ;
  RECT 353.460 0.000 354.580 1.120 ;
 END
END DI[20]
PIN DO[19]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal3 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal2 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal1 ;
  RECT 348.500 0.000 349.620 1.120 ;
 END
END DO[19]
PIN DI[19]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 340.440 0.000 341.560 1.120 ;
  LAYER metal3 ;
  RECT 340.440 0.000 341.560 1.120 ;
  LAYER metal2 ;
  RECT 340.440 0.000 341.560 1.120 ;
  LAYER metal1 ;
  RECT 340.440 0.000 341.560 1.120 ;
 END
END DI[19]
PIN DO[18]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal3 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal2 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal1 ;
  RECT 335.480 0.000 336.600 1.120 ;
 END
END DO[18]
PIN DI[18]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 326.800 0.000 327.920 1.120 ;
  LAYER metal3 ;
  RECT 326.800 0.000 327.920 1.120 ;
  LAYER metal2 ;
  RECT 326.800 0.000 327.920 1.120 ;
  LAYER metal1 ;
  RECT 326.800 0.000 327.920 1.120 ;
 END
END DI[18]
PIN DO[17]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 318.740 0.000 319.860 1.120 ;
  LAYER metal3 ;
  RECT 318.740 0.000 319.860 1.120 ;
  LAYER metal2 ;
  RECT 318.740 0.000 319.860 1.120 ;
  LAYER metal1 ;
  RECT 318.740 0.000 319.860 1.120 ;
 END
END DO[17]
PIN DI[17]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 310.060 0.000 311.180 1.120 ;
  LAYER metal3 ;
  RECT 310.060 0.000 311.180 1.120 ;
  LAYER metal2 ;
  RECT 310.060 0.000 311.180 1.120 ;
  LAYER metal1 ;
  RECT 310.060 0.000 311.180 1.120 ;
 END
END DI[17]
PIN DO[16]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 305.100 0.000 306.220 1.120 ;
  LAYER metal3 ;
  RECT 305.100 0.000 306.220 1.120 ;
  LAYER metal2 ;
  RECT 305.100 0.000 306.220 1.120 ;
  LAYER metal1 ;
  RECT 305.100 0.000 306.220 1.120 ;
 END
END DO[16]
PIN WEB[2]
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 300.760 0.000 301.880 1.120 ;
  LAYER metal3 ;
  RECT 300.760 0.000 301.880 1.120 ;
  LAYER metal2 ;
  RECT 300.760 0.000 301.880 1.120 ;
  LAYER metal1 ;
  RECT 300.760 0.000 301.880 1.120 ;
 END
END WEB[2]
PIN DI[16]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 297.040 0.000 298.160 1.120 ;
  LAYER metal3 ;
  RECT 297.040 0.000 298.160 1.120 ;
  LAYER metal2 ;
  RECT 297.040 0.000 298.160 1.120 ;
  LAYER metal1 ;
  RECT 297.040 0.000 298.160 1.120 ;
 END
END DI[16]
PIN A[1]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 290.840 0.000 291.960 1.120 ;
  LAYER metal3 ;
  RECT 290.840 0.000 291.960 1.120 ;
  LAYER metal2 ;
  RECT 290.840 0.000 291.960 1.120 ;
  LAYER metal1 ;
  RECT 290.840 0.000 291.960 1.120 ;
 END
END A[1]
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER metal4 ;
  RECT 284.640 0.000 285.760 1.120 ;
  LAYER metal3 ;
  RECT 284.640 0.000 285.760 1.120 ;
  LAYER metal2 ;
  RECT 284.640 0.000 285.760 1.120 ;
  LAYER metal1 ;
  RECT 284.640 0.000 285.760 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER metal4 ;
  RECT 282.780 0.000 283.900 1.120 ;
  LAYER metal3 ;
  RECT 282.780 0.000 283.900 1.120 ;
  LAYER metal2 ;
  RECT 282.780 0.000 283.900 1.120 ;
  LAYER metal1 ;
  RECT 282.780 0.000 283.900 1.120 ;
 END
END CS
PIN A[2]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 261.080 0.000 262.200 1.120 ;
  LAYER metal3 ;
  RECT 261.080 0.000 262.200 1.120 ;
  LAYER metal2 ;
  RECT 261.080 0.000 262.200 1.120 ;
  LAYER metal1 ;
  RECT 261.080 0.000 262.200 1.120 ;
 END
END A[2]
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER metal4 ;
  RECT 257.980 0.000 259.100 1.120 ;
  LAYER metal3 ;
  RECT 257.980 0.000 259.100 1.120 ;
  LAYER metal2 ;
  RECT 257.980 0.000 259.100 1.120 ;
  LAYER metal1 ;
  RECT 257.980 0.000 259.100 1.120 ;
 END
END CK
PIN A[0]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 256.120 0.000 257.240 1.120 ;
  LAYER metal3 ;
  RECT 256.120 0.000 257.240 1.120 ;
  LAYER metal2 ;
  RECT 256.120 0.000 257.240 1.120 ;
  LAYER metal1 ;
  RECT 256.120 0.000 257.240 1.120 ;
 END
END A[0]
PIN A[3]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER metal3 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER metal2 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER metal1 ;
  RECT 251.780 0.000 252.900 1.120 ;
 END
END A[3]
PIN A[4]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER metal3 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER metal2 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER metal1 ;
  RECT 244.340 0.000 245.460 1.120 ;
 END
END A[4]
PIN A[5]
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal3 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal2 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal1 ;
  RECT 241.240 0.000 242.360 1.120 ;
 END
END A[5]
PIN DO[15]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal3 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal2 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal1 ;
  RECT 233.180 0.000 234.300 1.120 ;
 END
END DO[15]
PIN DI[15]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal3 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal2 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal1 ;
  RECT 224.500 0.000 225.620 1.120 ;
 END
END DI[15]
PIN DO[14]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal3 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal2 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal1 ;
  RECT 219.540 0.000 220.660 1.120 ;
 END
END DO[14]
PIN DI[14]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal3 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal2 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal1 ;
  RECT 211.480 0.000 212.600 1.120 ;
 END
END DI[14]
PIN DO[13]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal3 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal2 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal1 ;
  RECT 202.800 0.000 203.920 1.120 ;
 END
END DO[13]
PIN DI[13]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal3 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal2 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal1 ;
  RECT 194.740 0.000 195.860 1.120 ;
 END
END DI[13]
PIN DO[12]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal3 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal2 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal1 ;
  RECT 189.780 0.000 190.900 1.120 ;
 END
END DO[12]
PIN DI[12]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal3 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal2 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal1 ;
  RECT 181.100 0.000 182.220 1.120 ;
 END
END DI[12]
PIN DO[11]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal3 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal2 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal1 ;
  RECT 176.140 0.000 177.260 1.120 ;
 END
END DO[11]
PIN DI[11]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal3 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal2 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal1 ;
  RECT 168.080 0.000 169.200 1.120 ;
 END
END DI[11]
PIN DO[10]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal3 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal2 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal1 ;
  RECT 163.120 0.000 164.240 1.120 ;
 END
END DO[10]
PIN DI[10]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal3 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal2 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal1 ;
  RECT 154.440 0.000 155.560 1.120 ;
 END
END DI[10]
PIN DO[9]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO[9]
PIN DI[9]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal3 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal2 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal1 ;
  RECT 137.700 0.000 138.820 1.120 ;
 END
END DI[9]
PIN DO[8]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO[8]
PIN WEB[1]
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 128.400 0.000 129.520 1.120 ;
  LAYER metal3 ;
  RECT 128.400 0.000 129.520 1.120 ;
  LAYER metal2 ;
  RECT 128.400 0.000 129.520 1.120 ;
  LAYER metal1 ;
  RECT 128.400 0.000 129.520 1.120 ;
 END
END WEB[1]
PIN DI[8]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI[8]
PIN DO[7]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO[7]
PIN DI[7]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI[7]
PIN DO[6]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO[6]
PIN DI[6]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI[6]
PIN DO[5]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO[5]
PIN DI[5]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI[5]
PIN DO[4]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO[4]
PIN DI[4]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI[4]
PIN DO[3]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO[3]
PIN DI[3]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI[3]
PIN DO[2]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO[2]
PIN DI[2]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI[2]
PIN DO[1]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO[1]
PIN DI[1]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI[1]
PIN DO[0]
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO[0]
PIN WEB[0]
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 15.560 0.000 16.680 1.120 ;
  LAYER metal3 ;
  RECT 15.560 0.000 16.680 1.120 ;
  LAYER metal2 ;
  RECT 15.560 0.000 16.680 1.120 ;
  LAYER metal1 ;
  RECT 15.560 0.000 16.680 1.120 ;
 END
END WEB[0]
PIN DI[0]
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI[0]
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 531.960 156.800 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 531.960 156.800 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 531.960 156.800 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 531.960 156.800 ;
  LAYER via ;
  RECT 0.000 0.140 531.960 156.800 ;
  LAYER via2 ;
  RECT 0.000 0.140 531.960 156.800 ;
  LAYER via3 ;
  RECT 0.000 0.140 531.960 156.800 ;
END
END data_array
END LIBRARY



